module test6(a,b);
input [7:0]a;
output [7:0]b;
wire [7:0]a,b;
assign b=a;
endmodule 